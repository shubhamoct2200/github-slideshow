//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Assignment5.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w16;    //: /sn:0 {0}(91,207)(101,207)(101,158)(121,158){1}
supply0 w0;    //: /sn:0 {0}(462,176)(462,194)(412,194)(412,209){1}
reg [7:0] w3;    //: /sn:0 {0}(#:235,527)(266,527)(266,388){1}
//: {2}(266,384)(266,308)(274,308){3}
//: {4}(278,308)(339,308){5}
//: {6}(343,308)(355,308){7}
//: {8}(#:359,308)(516,308)(516,350){9}
//: {10}(357,310)(357,341){11}
//: {12}(341,306)(341,163)(346,163)(346,153){13}
//: {14}(348,151)(444,151){15}
//: {16}(344,151)(321,151)(#:321,130){17}
//: {18}(276,306)(276,274)(#:204,274){19}
//: {20}(264,386)(245,386)(245,385)(#:203,385){21}
reg w20;    //: /sn:0 {0}(98,443)(116,443)(116,449)(129,449){1}
reg w29;    //: /sn:0 {0}(454,451)(464,451)(464,478)(407,478)(407,498){1}
reg w19;    //: /sn:0 {0}(195,380)(195,372)(234,372)(234,357)(229,357){1}
reg w18;    //: /sn:0 {0}(96,317)(103,317)(103,312)(113,312){1}
reg w21;    //: /sn:0 {0}(230,490)(239,490)(239,514)(227,514)(227,522){1}
reg w17;    //: /sn:0 {0}(196,269)(196,250)(207,250)(207,235)(197,235){1}
reg w27;    //: /sn:0 {0}(566,321)(582,321)(582,364)(524,364){1}
reg w28;    //: /sn:0 {0}(556,410)(556,373)(664,373)(664,411)(636,411){1}
supply0 w2;    //: /sn:0 {0}(229,415)(229,413){1}
//: {2}(229,409)(229,347){3}
//: {4}(229,343)(229,163)(197,163){5}
//: {6}(227,345)(196,345)(196,317)(189,317){7}
//: {8}(227,411)(210,411)(210,454)(205,454){9}
reg w15;    //: /sn:0 {0}(205,444)(237,444)(237,338){1}
//: {2}(237,334)(237,296)(234,296)(234,262){3}
//: {4}(234,258)(234,100)(204,100){5}
//: {6}(232,260)(212,260)(212,153)(197,153){7}
//: {8}(235,336)(202,336)(202,307)(189,307){9}
wire [7:0] w6;    //: /sn:0 {0}(#:134,249)(134,274)(156,274){1}
//: {2}(160,274)(188,274){3}
//: {4}(#:158,272)(#:158,169){5}
wire [7:0] w13;    //: /sn:0 {0}(#:308,387)(308,411)(370,411){1}
//: {2}(374,411)(383,411)(383,382)(373,382)(#:373,370){3}
//: {4}(#:372,413)(372,503)(399,503){5}
wire [7:0] w4;    //: /sn:0 {0}(#:415,503)(434,503)(434,597){1}
//: {2}(436,599)(567,599)(567,415)(#:564,415){3}
//: {4}(432,599)(320,599){5}
//: {6}(318,597)(318,595)(319,595)(#:319,561){7}
//: {8}(316,599)(46,599)(46,401){9}
//: {10}(48,399)(166,399)(#:166,439){11}
//: {12}(46,397)(46,288){13}
//: {14}(#:48,286)(150,286)(150,302){15}
//: {16}(46,284)(46,130)(158,130)(#:158,148){17}
wire [7:0] w10;    //: /sn:0 {0}(#:129,514)(129,527)(165,527){1}
//: {2}(169,527)(219,527){3}
//: {4}(#:167,525)(167,503)(166,503)(#:166,460){5}
wire [7:0] w24;    //: /sn:0 {0}(#:455,387)(455,415)(502,415){1}
//: {2}(506,415)(548,415){3}
//: {4}(#:504,413)(504,409)(500,409)(#:500,379){5}
wire [7:0] w1;    //: /sn:0 {0}(589,124)(589,149)(#:479,149){1}
wire [7:0] w11;    //: /sn:0 {0}(#:389,341)(389,322)(#:484,322)(484,350){1}
wire [7:0] w5;    //: /sn:0 {0}(#:89,370)(89,375)(171,375){1}
//: {2}(173,373)(173,339)(150,339)(#:150,323){3}
//: {4}(173,377)(173,385)(187,385){5}
wire w26;    //: /sn:0 {0}(452,345)(452,364)(476,364){1}
//: enddecls

  //: comment g8 @(446,115) /sn:0
  //: /line:"ROM"
  //: /end
  //: frame g4 @(247,82) /sn:0 /wi:426 /ht:151 /tx:""
  //: GROUND g3 (w0) @(412,215) /sn:0 /w:[ 1 ]
  //: SWITCH g16 (w28) @(619,411) /sn:0 /w:[ 1 ] /st:1 /dn:1
  //: joint g47 (w4) @(318, 599) /w:[ 5 6 8 -1 ]
  //: joint g26 (w3) @(266, 386) /w:[ -1 2 20 1 ]
  //: SWITCH g17 (w29) @(437,451) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g2 (w1) @(589,117) /sn:0 /w:[ 0 ] /type:1
  //: joint g30 (w5) @(173, 375) /w:[ -1 2 1 4 ]
  //: LED g23 (w10) @(129,507) /sn:0 /w:[ 0 ] /type:1
  //: joint g39 (w3) @(341, 308) /w:[ 6 12 5 -1 ]
  //: DIP g1 (w3) @(321,120) /sn:0 /w:[ 17 ] /st:2 /dn:1
  //: LED g24 (w5) @(89,363) /sn:0 /w:[ 0 ] /type:1
  //: joint g29 (w3) @(276, 308) /w:[ 4 18 3 -1 ]
  _GGBUFIF8 #(4, 6) g51 (.Z(w3), .I(w5), .E(w19));   //: @(193,385) /sn:0 /w:[ 21 5 0 ]
  //: joint g18 (w13) @(372, 411) /w:[ 2 -1 1 4 ]
  //: SWITCH g10 (w20) @(81,443) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g25 (w6) @(134,242) /sn:0 /w:[ 0 ] /type:1
  //: joint g49 (w2) @(229, 345) /w:[ -1 4 6 3 ]
  //: comment g6 @(569,92) /sn:0
  //: /line:"led bar"
  //: /end
  _GGBUFIF8 #(4, 6) g50 (.Z(w3), .I(w6), .E(w17));   //: @(194,274) /sn:0 /w:[ 19 3 0 ]
  //: comment g9 @(254,71) /sn:0
  //: /line:"ROM INPUT"
  //: /end
  //: comment g7 @(288,86) /sn:0
  //: /line:"DIP Switch"
  //: /end
  //: LED g35 (w26) @(452,338) /sn:0 /w:[ 0 ] /type:0
  //: joint g56 (w4) @(434, 599) /w:[ 2 1 4 -1 ]
  _GGMUL8 #(124) g58 (.A(w3), .B(w11), .P(w13));   //: @(373,357) /sn:0 /w:[ 11 0 3 ]
  //: LED g22 (w4) @(319,554) /sn:0 /w:[ 7 ] /type:1
  //: joint g31 (w4) @(46, 286) /w:[ 14 16 -1 13 ]
  //: joint g33 (w15) @(237, 336) /w:[ -1 2 8 1 ]
  //: joint g36 (w2) @(229, 411) /w:[ -1 2 8 1 ]
  _GGBUFIF8 #(4, 6) g41 (.Z(w4), .I(w24), .E(w28));   //: @(554,415) /sn:0 /w:[ 3 3 0 ]
  //: joint g42 (w3) @(346, 151) /w:[ 14 -1 16 13 ]
  _GGBUFIF8 #(4, 6) g52 (.Z(w3), .I(w10), .E(w21));   //: @(225,527) /sn:0 /w:[ 0 3 1 ]
  //: joint g40 (w3) @(357, 308) /w:[ 8 -1 7 10 ]
  _GGREG8 #(10, 10, 20) g12 (.Q(w10), .D(w4), .EN(w2), .CLR(w15), .CK(w20));   //: @(166,449) /sn:0 /w:[ 5 11 9 0 1 ]
  _GGBUFIF8 #(4, 6) g34 (.Z(w4), .I(w13), .E(w29));   //: @(405,503) /sn:0 /w:[ 0 5 1 ]
  //: joint g28 (w6) @(158, 274) /w:[ 2 4 1 -1 ]
  //: joint g46 (w4) @(46, 399) /w:[ 10 12 -1 9 ]
  //: SWITCH g5 (w16) @(74,207) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g11 (w15) @(187,100) /sn:0 /w:[ 5 ] /st:1 /dn:1
  //: GROUND g14 (w2) @(229,421) /sn:0 /w:[ 0 ]
  //: SWITCH g19 (w19) @(212,357) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: joint g21 (w15) @(234, 260) /w:[ -1 4 6 3 ]
  //: SWITCH g20 (w21) @(213,490) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGADD8 #(68, 70, 62, 64) g32 (.A(w11), .B(w3), .S(w24), .CI(w27), .CO(w26));   //: @(500,366) /sn:0 /w:[ 1 9 5 1 1 ]
  _GGROM8x8 #(10, 30) g0 (.A(w3), .D(w1), .OE(w0));   //: @(462,150) /sn:0 /w:[ 15 1 0 ] /mem:"/home/sam/Downloads/test.mem"
  //: SWITCH g15 (w18) @(79,317) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: LED g38 (w13) @(308,380) /sn:0 /w:[ 0 ] /type:1
  //: LED g43 (w24) @(455,380) /sn:0 /w:[ 0 ] /type:1
  //: SWITCH g27 (w17) @(180,235) /sn:0 /w:[ 1 ] /st:1 /dn:1
  _GGREG8 #(10, 10, 20) g48 (.Q(w5), .D(w4), .EN(w2), .CLR(w15), .CK(w18));   //: @(150,312) /sn:0 /w:[ 3 15 7 9 1 ]
  //: joint g37 (w24) @(504, 415) /w:[ 2 4 1 -1 ]
  //: joint g55 (w10) @(167, 527) /w:[ 2 4 1 -1 ]
  _GGREG8 #(10, 10, 20) g13 (.Q(w6), .D(w4), .EN(w2), .CLR(w15), .CK(w16));   //: @(158,158) /sn:0 /w:[ 5 17 5 7 1 ]
  //: SWITCH g53 (w27) @(549,321) /sn:0 /w:[ 0 ] /st:0 /dn:1

endmodule
//: /netlistEnd

